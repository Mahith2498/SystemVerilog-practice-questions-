`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Create Date: 02/07/2026 12:59:14 PM
// Designer Name: KOTHAPALLI MAHITH VATHSAV 
// Module Name: tbone
// Project Name: Hello SystemVerilog program  
module tbone;
string prog = "Hello SystemVerilog!!";
initial begin 
$display("%s",prog);
end
endmodule
